
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:29:09 11/18/2022 
// Design Name: 
// Module Name:    Timer0 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
`define IDLE 2'b00
`define LOAD 2'b01
`define CNT  2'b10
`define INT  2'b11

`define ctrl   mem[0]
`define preset mem[1]
`define count  mem[2]
module Timer(
    input clk,
    input reset,
    input [31:0] Addr,
    input WE,
    input [31:0] Din,
    output [31:0] Dout,
    output IRQ
    );

	reg [1:0] state;
	reg [31:0] mem [2:0];
	
	reg _IRQ;
	assign IRQ = `ctrl[3] & _IRQ;
	
	assign Dout = mem[Addr[3:2]];
	
	wire [31:0] load = Addr[3:2] == 2'b0 ? {28'h0, Din[3:0]} : Din;
	
	localparam PERIOD = 32'd25000000; // clk is 25MHz
	reg [31:0] counter;
    always @(posedge clk) begin
        if (reset) 
            counter <= 0;
        else begin
            if (counter + 1 == PERIOD || state == `IDLE)
                counter <= 0;
            else
                counter <= counter + 1;
        end
    end
	integer i;
	always @(posedge clk) begin
		if(reset) begin
			state <= 0; 
			for(i = 0; i < 3; i = i+1) mem[i] <= 0;
			_IRQ <= 0;
		end
		else if(WE) begin
			// $display("%d@: *%h <= %h", $time, {Addr, 2'b00}, load);
			mem[Addr[3:2]] <= load;
		end
		if (reset != 1) begin
			case(state)
				`IDLE : if(`ctrl[0]) begin
					state <= `LOAD;
					_IRQ <= 1'b0;
				end
				`LOAD : begin
					if(`ctrl[2:1] == 2'b00 || `ctrl[2:1] == 2'b01) begin
							`count <= `preset;
					end
					else if(`ctrl[2:1] == 2'b10) begin
							`count <= 0;
					end
					state <= `CNT;
				end
				`CNT  : 
					if(WE == 1 & Din != `preset & Addr[3:2] == 1) begin
							state <= `IDLE;
					end
					else if(`ctrl[0]) begin
						if(`count > 1 && counter + 1 == PERIOD && (`ctrl[2:1] == 2'b00 || `ctrl[2:1] == 2'b01)) begin 
								`count <= `count-1;
						end
						else if(`count < `preset -1 && counter + 1 == PERIOD && `ctrl[2:1] == 2'b10) begin
								`count <= `count + 1;
						end
						else if (`count == 1 && counter + 1 == PERIOD && (`ctrl[2:1] == 2'b00 || `ctrl[2:1] == 2'b01)) begin
							`count <= 0;
							state <= `INT;
							_IRQ <= 1'b1;
						end
						else if (`count == `preset - 1 && counter + 1 == PERIOD && `ctrl[2:1] == 2'b10) begin
							`count <= `preset;
							state <= `INT;
							_IRQ <= 1'b1;
						end
						else if(`preset == 0 && `ctrl[2:1] == 2'b10) begin
							`count <= 0;
							state <= `INT;
							_IRQ <= 1'b1;
						end
					end
					else state <= `IDLE;
				default : begin
					if(counter + 1 == PERIOD) begin
						if(`ctrl[2:1] == 2'b00 || `ctrl[2:1] == 2'b10) `ctrl[0] <= 1'b0;
						else _IRQ <= 1'b0;
						state <= `IDLE;
					end
				end
			endcase
		end
	end

endmodule

