`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:45:30 12/06/2022 
// Design Name: 
// Module Name:    M_RegDstSel 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module M_RegDstSel(
    input [4:0] M_A3,
    input [4:0] M_A3FromDM,
    output [4:0] M_TrueA3,
    input M_Check
    );


endmodule
